package uvmtb_sequence_pkg;
	import uvm_pkg::*;
	import uvmtb_keypad_agent_pkg::Alu_packet;
	import uvmtb_keypad_agent_pkg::Key;
	import utils_pkg::*;
	`include "uvm_macros.svh"
	`include "uvmtb_sequence_random.svh"
	`include "uvmtb_sequence_2ndOperand_equal_0.svh"
	`include "uvmtb_sequence_single_digit_operation.svh"
	`include "uvmtb_virtual_sequence.svh"

endpackage