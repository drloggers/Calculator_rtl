package uvmtb_display_agent_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "Result.svh"
	import uvmtb_keypad_agent_pkg::*;
	import utils_pkg::*;
	`include "uvmtb_display_config.svh"
	`include "uvmtb_display_driver.svh"
	`include "uvmtb_display_monitor.svh"
	`include "uvmtb_display_key_monitor.svh"
	`include "uvmtb_display_agent.svh"
endpackage