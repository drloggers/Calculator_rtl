package utils_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	`include "utils_functions.svh"

endpackage